`timescale 1ns/1ps
`include "ALU.v"

module alu_test;

reg[31:0] instruction, regA, regB;

wire[31:0] result;
wire[2:0] flags;

alu testalu(instruction, regA, regB, result, flags);

initial
begin

$dumpfile("test_ALU.vcd");
$dumpvars(0, alu_test);

$display("Format of output");
$monitor("instruction\t= %32b \nop\t\t= %6b \nfunc\t\t= %6b \nreg_A\t\t= %h \nreg_B\t\t= %h \nreg_rs\t\t= %h \nreg_regB\t\t= %h \nresult\t\t= %h \nflags\t\t= %3b \n",
instruction, test_alu.opcode, test_alu.func, regA, regB, test_alu.rs, test_alu.rt, result, flags);

// 1. add
#10 instruction<=32'b0000_0000_0000_0001_0110_0000_0010_0000;   //add $t4, regA, regB
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0000; 


// 2. addi
#10 instruction<=32'b0010_0000_0000_1111_0000_0000_0000_1010;   //addi $t7, regA, 10
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0110;

// 3. addu
#10 instruction<=32'b0000_0000_0000_0001_0110_0000_0010_0001;   //addu $t4, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_0010;

// 4. addiu
#10 instruction<=32'b0010_0100_0000_1111_0000_0000_0000_1010;   //addiu $t7, regA, 10
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0110;

// 5. sub
#10 instruction <= 32'b0000_0000_0000_0001_0000_1000_0010_0010; //sub $at, $reg_A, $reg_B
regA <= 32'b1111_1111_1111_1111_1111_1111_1101_1101;
regB <= 32'b0000_0000_0000_0000_0000_0000_0010_0101;

// 6. subu
#10 instruction<=32'b0000_0000_0000_0001_0100_0000_0010_0011;   //subu $t0, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_0001_0010;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_1010;

// 7. and
#10 instruction<=32'b0000_0000_0000_0001_0110_1000_0010_0100;   //and $t5, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_1101;

// 8. andi
#10 instruction<=32'b0011_0000_0000_1101_0000_0000_0000_1001;   //and $t5, regA, 9
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

// 9. nor
#10 instruction<=32'b0000_0000_0000_0001_0111_0000_0010_0111;   //nor $t6, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_1101;

// 10. or
#10 instruction<=32'b0000_0000_0000_0001_0111_0000_0010_0101;   //or $t6, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_1001_0110;
regB<=32'b0000_0000_0000_0000_0000_0100_1101_1101;

// 11. ori
#10 instruction<=32'b0011_0100_0000_1010_1111_1111_1111_0001;   //ori $t2, regA, -15
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

// 12. xor
#10 instruction<=32'b0000_0000_0000_0001_0111_0000_0010_0110;   //xor $t6, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
regB<=32'b0000_0000_0000_0000_0000_0100_1101_1101;

// 13. xori
#10 instruction<=32'b0011_1000_0000_1010_1111_1111_1111_0001;   //xori $t2, regA, -15
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

// 14. beq
#10 instruction<=32'b0001_0000_0010_0000_0000_0000_0000_1010;   //beq regA, regB, 10
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

// 15. bne
#10 instruction<=32'b0001_0100_0000_0001_0000_0000_0000_0111;   //bne regA, regB, 7
regA<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

// 16. slt
#10 instruction<=32'b0000_0000_0000_0001_0111_1000_0010_1010;   //slt $t1, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

// 17. slti
#10 instruction<=32'b0010_1000_0001_0001_0000_0000_0000_1101;   //slti $s1, regA, 13
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

// 18. sltiu
#10 instruction<=32'b0010_1100_0001_0001_1111_1111_1111_0011;   //sltiu $s1, regA, -13
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

// 19. sltu
#10 instruction<=32'b0000_0000_0000_0001_0111_1000_0010_1011;   //sltu $t1, regA, regB
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_1000;

// 20. lw
#10 instruction <= 32'b1000_1100_0011_0000_0000_0000_0000_0000; //lw $s0, 0($regB)
regB <= 32'b0000_0000_0000_0000_0000_1000_0001_0000;

// 21. sw
#10 instruction <= 32'b1010_1100_0000_1001_0000_0000_0000_1010; //sw $t1, 10($reg_A)
reg_A <= 32'b0000_0000_0000_0000_0000_0000_1100_0100;

// 22. sll
#10 instruction<=32'b0000_0000_0000_0001_0110_0001_0100_0000;   //sll $t4, regB, 5
regB<=32'b1001_1001_1111_1111_1001_1001_1101_1101;

// 23. sllv
#10 instruction<=32'b0000_0000_0000_0001_0110_0000_0000_0100;   //sllv $t4, regB, regA
regB<=32'b1001_1001_1111_1111_1001_1001_1101_1101;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

// 24. srl
#10 instruction<=32'b0000_0000_0000_0001_0110_0001_0100_0010;   //srl $t4, regB, 5
regB<=32'b1001_1001_1111_1111_1001_1001_1101_1101;

// 25. srlv
#10 instruction<=32'b0000_0000_0000_0001_0110_0000_0000_0110;   //srlv $t4, regB, regA
regB<=32'b1001_1001_1111_1111_1001_1001_1101_1101;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

// 26. sra
#10 instruction <= 32'b0000_0000_0010_0000_0111_1000_1000_0011; //sra $t5, $reg_A, 2
reg_A <= 32'b1001_1001_1111_1111_1001_1001_1101_1101;

// 27. srav
#10 instruction <= 32'b0000_0000_0010_0000_1100_0000_0000_0111; //srav $t8, $reg_A, $reg_B
reg_A <= 32'b1001_1001_1111_1111_1001_1001_1101_1101;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;


#10 $finish;
end
endmodule